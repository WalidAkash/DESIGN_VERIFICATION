// Description here
// ### Author : name (email)

module tb_reg_file;

  //`define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "../include/tb_ess.sv"

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  localparam int ADW = 5;
  localparam int DPW = 32;



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:3 tLow:7
  `CREATE_CLK(clk_i, 3, 7)
  logic [ADW-1:0] addr_1;
  logic [ADW-1:0] addr_2;
  logic [ADW-1:0] addr_3;
  logic           we;
  logic [DPW-1:0] wd_3;
  logic [DPW-1:0] rd_1;
  logic [DPW-1:0] rd_2;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////
  logic [DPW-1:0] regs_mem[0:((2**ADW)-1)];


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  /* assign regs[addr_1] = [DPW-1:0]regs_mem[0];
  assign regs[addr_2] = [DPW-1:0]regs_mem[1];
  assign regs[addr_3] = [DPW-1:0]regs_mem[2]; */


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////
  reg_file #(
    .ADW(ADW),
    .DPW(DPW)
) dut (
    .clk_i(clk_i),
    .addr_1(addr_1),
    .addr_2(addr_2),
    .addr_3(addr_3),
    .we(we),
    .wd_3(wd_3),
    .rd_1(rd_1),
    .rd_2(rd_2)
);


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin
    start_clk_i();
    @(posedge clk_i);


    /*
    // Write data to addr_3
    addr_3 = 2;
    we = 1;
    wd_3 = 32'h12345678;
    #10;
    we = 0;

    // Read data from addr_1 and addr_2
    addr_1 = 0;
    addr_2 = 1;
    #10;

    // Verify results
    if (rd_1 !== 32'h00000000) $error("Test failed: rd_1");
    if (rd_2 !== 32'h00000000) $error("Test failed: rd_2");

    addr_1 = 2;
    addr_2 = 2;
    #10;

    if (rd_1 !== 32'h12345678) $error("Test failed: rd_1");
    if (rd_2 !== 32'h12345678) $error("Test failed: rd_2");*/

    $display("Test passed");
    #100;
    $finish;
  end

endmodule
