// Designer : Walid Akash
// Company : DSi
// Description : decode stage pipeline register

module top_stage
  import rv32i_pkg::*;
();

endmodule
