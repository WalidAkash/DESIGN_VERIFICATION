module riscv(
  
);

endmodule