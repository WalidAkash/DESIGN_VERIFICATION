// Designer : Walid Akash
// Company : DSi

module tb_decode_stage;
import rv32i_pkg::*;


endmodule