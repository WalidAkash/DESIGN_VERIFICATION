// Designer : Walid Akash
// Company : DSi
// Description : This module shifts the instruction by an appropriate amount

module extend_unit (
    input  logic [31:7] instr,
    input  logic [ 1:0] immsrc,
    output logic [31:0] immext
);



endmodule
