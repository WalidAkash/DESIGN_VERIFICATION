// Designer : Walid Akash
// Company : DSi

module branch_unit;

endmodule